library verilog;
use verilog.vl_types.all;
entity Tb_filter_IIR is
    generic(
        Nb              : integer := 10
    );
end Tb_filter_IIR;
